// Global nets module 
`timescale 1ns / 1ns

`celldefine
module cds_globals;


supply1 vdd_;

supply0 gnd_;


endmodule
`endcelldefine
